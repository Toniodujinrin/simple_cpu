module simple_cpu(); 


endmodule 