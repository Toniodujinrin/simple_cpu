module hazard_detector()


endmodule 