module branch_controler(); 



endmodule 