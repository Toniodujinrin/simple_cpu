
//4-way set associative cache with write-back, write-allocate policy 

module cache(); 


endmodule