///////////////////////////////////////////////////////////////////////////////
// File:        ID_EX_reg.v
// Author:      Toni Odujinrin
// Date:        2025-10-04 
// Description: MEM_WB pipeline register 
///////////////////////////////////////////////////////////////////////////////


module MEM_WB_REG(


); 


endmodule 